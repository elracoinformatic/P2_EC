//: version "1.8.7"

module Shift_Left_2(out, in);
//: interface  /sz:(142, 98) /bd:[ Li0>in[25:0](42/98) Ro0<out[27:0](52/98) ]
input [25:0] in;    //: /sn:0 {0}(102,173)(290,173)(290,174)(300,174){1}
output [27:0] out;    //: /sn:0 {0}(424,216)(343,216)(343,184)(306,184){1}
supply0 w2;    //: /sn:0 {0}(182,248)(182,196){1}
//: {2}(184,194)(300,194){3}
//: {4}(182,192)(182,184)(300,184){5}
//: enddecls

  //: joint g4 (w2) @(182, 194) /w:[ 2 4 -1 1 ]
  //: supply0 g3 (w2) @(182,254) /sn:0 /w:[ 0 ]
  concat g2 (.I0(w2), .I1(w2), .I2(in), .Z(out));   //: @(305,184) /sn:0 /w:[ 3 5 1 1 ] /dr:0
  //: output g1 (out) @(421,216) /sn:0 /w:[ 0 ]
  //: input g0 (in) @(100,173) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [25:0] w0;    //: /sn:0 {0}(213,115)(223,115){1}
wire [27:0] w1;    //: /sn:0 {0}(377,125)(367,125){1}
//: enddecls

  Shift_Left_2 g0 (.in(w0), .out(w1));   //: @(224, 73) /sz:(142, 98) /sn:0 /p:[ Li0>1 Ro0<1 ]

endmodule
