//: version "1.8.7"

module EXE(ALU_result, Zero, B, A, ALU_operation);
//: interface  /sz:(182, 314) /bd:[ Ti0>ALU_operation[3:0](84/182) Li0>B[31:0](132/314) Li1>A[31:0](66/314) Ro0<Zero(65/314) Ro1<ALU_result[31:0](135/314) ]
input [31:0] B;    //: /sn:0 {0}(166,377)(387,377){1}
output Zero;    //: /sn:0 {0}(540,308)(675,308){1}
output [31:0] ALU_result;    //: /sn:0 {0}(540,374)(679,374){1}
input [31:0] A;    //: /sn:0 {0}(170,301)(387,301){1}
input [3:0] ALU_operation;    //: /sn:0 {0}(406,120)(464,120)(464,244){1}
//: enddecls

  //: output g4 (ALU_result) @(676,374) /sn:0 /w:[ 1 ]
  //: output g3 (Zero) @(672,308) /sn:0 /w:[ 1 ]
  //: input g2 (B) @(164,377) /sn:0 /w:[ 0 ]
  //: input g1 (A) @(168,301) /sn:0 /w:[ 0 ]
  //: input g5 (ALU_operation) @(404,120) /sn:0 /w:[ 0 ]
  ALU g0 (.ALU_operation(ALU_operation), .B(B), .A(A), .ALU_result(ALU_result), .Zero(Zero));   //: @(388, 245) /sz:(151, 203) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<0 Ro1<0 ]

endmodule

module ALU(B, ALU_operation, ALU_result, A, Zero);
//: interface  /sz:(127, 166) /bd:[ Ti0>ALU_operation[3:0](64/127) Li0>B[31:0](108/166) Li1>A[31:0](46/166) Ro0<ALU_result[31:0](106/166) Ro1<Zero(52/166) ]
supply0 w7;    //: /sn:0 /dp:1 {0}(651,129)(651,110){1}
input [31:0] B;    //: /sn:0 {0}(415,270)(468,270){1}
//: {2}(472,270)(594,270){3}
//: {4}(598,270)(643,270){5}
//: {6}(647,270)(700,270)(700,302)(743,302){7}
//: {8}(645,272)(645,370)(720,370){9}
//: {10}(596,272)(596,392)(718,392){11}
//: {12}(470,268)(470,207)(471,207){13}
output Zero;    //: /sn:0 /dp:1 {0}(1222,354)(1270,354){1}
output [31:0] ALU_result;    //: /sn:0 /dp:1 {0}(1029,324)(1134,324)(1134,322)(1144,322){1}
//: {2}(1146,320)(1146,292)(1194,292){3}
//: {4}(1146,324)(1146,351)(1201,351){5}
supply0 w3;    //: /sn:0 /dp:1 {0}(552,145)(552,123){1}
supply0 w0;    //: /sn:0 {0}(757,243)(757,262){1}
input [31:0] A;    //: /sn:0 {0}(412,238)(610,238){1}
//: {2}(614,238)(659,238){3}
//: {4}(663,238)(708,238)(708,270)(743,270){5}
//: {6}(661,240)(661,365)(720,365){7}
//: {8}(612,236)(612,137)(637,137){9}
//: {10}(612,240)(612,387)(718,387){11}
supply0 [31:0] w20;    //: /sn:0 {0}(805,115)(805,119)(899,119){1}
input [3:0] ALU_operation;    //: /sn:0 {0}(428,544)(722,544)(722,543)(1015,543){1}
//: {2}(1016,543)(1077,543){3}
supply0 [31:0] w1;    //: /sn:0 {0}(1166,382)(1166,369)(1185,369)(1185,359){1}
//: {2}(1187,357)(1188,357)(1188,356)(1201,356){3}
//: {4}(1183,357)(1178,357){5}
supply0 [31:0] w5;    //: /sn:0 {0}(825,318)(857,318)(857,317)(867,317){1}
//: {2}(869,315)(869,314)(1000,314){3}
//: {4}(869,319)(869,320)(983,320){5}
//: {6}(987,320)(1000,320){7}
//: {8}(985,322)(985,327)(1000,327){9}
wire [31:0] w16;    //: /sn:0 {0}(666,153)(818,153)(818,159){1}
//: {2}(818,160)(818,307)(1000,307){3}
wire [31:0] w6;    //: /sn:0 {0}(567,169)(637,169){1}
wire w4;    //: /sn:0 {0}(757,310)(757,338){1}
wire w19;    //: /sn:0 {0}(651,177)(651,197){1}
wire [31:0] w12;    //: /sn:0 {0}(487,207)(512,207)(512,185)(538,185){1}
wire [31:0] w18;    //: /sn:0 {0}(741,368)(793,368)(793,347)(1000,347){1}
wire [2:0] w10;    //: /sn:0 {0}(1016,538)(1016,347){1}
wire w8;    //: /sn:0 {0}(552,193)(552,203)(565,203)(565,213){1}
wire [31:0] w17;    //: /sn:0 {0}(928,109)(990,109)(990,300)(1000,300){1}
wire [31:0] w11;    //: /sn:0 {0}(465,133)(465,153)(518,153){1}
//: {2}(522,153)(538,153){3}
//: {4}(520,151)(520,99)(899,99){5}
wire [31:0] w2;    //: /sn:0 {0}(772,286)(800,286)(800,334)(1000,334){1}
wire w15;    //: /sn:0 {0}(822,160)(915,160)(915,132){1}
wire [31:0] w9;    //: /sn:0 {0}(739,390)(803,390)(803,340)(1000,340){1}
//: enddecls

  //: joint g8 (A) @(612, 238) /w:[ 2 8 1 10 ]
  or g4 (.I0(A), .I1(B), .Z(w9));   //: @(729,390) /sn:0 /w:[ 11 11 0 ]
  //: supply0 g16 (w5) @(819,318) /sn:0 /R:3 /w:[ 0 ]
  and g3 (.I0(A), .I1(B), .Z(w18));   //: @(731,368) /sn:0 /w:[ 7 9 0 ]
  add g26 (.A(w6), .B(A), .S(w16), .CI(w7), .CO(w19));   //: @(653,153) /sn:0 /R:1 /w:[ 1 9 0 0 0 ]
  //: supply0 g17 (w1) @(1166,388) /sn:0 /w:[ 0 ]
  //: joint g2 (ALU_result) @(1146, 322) /w:[ -1 2 1 4 ]
  //: joint g30 (w5) @(869, 317) /w:[ -1 2 1 4 ]
  //: joint g23 (B) @(470, 270) /w:[ 2 12 1 -1 ]
  //: supply0 g24 (w3) @(552,117) /sn:0 /R:2 /w:[ 1 ]
  //: joint g1 (A) @(661, 238) /w:[ 4 -1 3 6 ]
  mux g29 (.I0(w18), .I1(w9), .I2(w2), .I3(w5), .I4(w5), .I5(w5), .I6(w16), .I7(w17), .S(w10), .Z(ALU_result));   //: @(1016,324) /sn:0 /R:1 /w:[ 1 1 1 9 7 3 3 1 1 0 ] /ss:0 /do:0
  //: joint g18 (w1) @(1185, 357) /w:[ 2 -1 4 1 ]
  led g25 (.I(w8));   //: @(565,220) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: supply0 g10 (w0) @(757,237) /sn:0 /R:2 /w:[ 0 ]
  //: input g6 (B) @(413,270) /sn:0 /w:[ 0 ]
  //: joint g35 (w11) @(520, 153) /w:[ 2 4 1 -1 ]
  //: joint g9 (B) @(596, 270) /w:[ 4 -1 3 10 ]
  //: joint g7 (B) @(645, 270) /w:[ 6 -1 5 8 ]
  //: joint g31 (w5) @(985, 320) /w:[ 6 -1 5 8 ]
  add g22 (.A(w12), .B(w11), .S(w6), .CI(w3), .CO(w8));   //: @(554,169) /sn:0 /R:1 /w:[ 1 3 0 0 0 ]
  tran g33(.Z(w15), .I(w16[31]));   //: @(816,160) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: input g12 (ALU_operation) @(426,544) /sn:0 /w:[ 0 ]
  //: supply0 g34 (w20) @(805,109) /sn:0 /R:2 /w:[ 0 ]
  led g28 (.I(w19));   //: @(651,204) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: output g14 (ALU_result) @(1191,292) /sn:0 /w:[ 3 ]
  led g11 (.I(w4));   //: @(757,345) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: input g5 (A) @(410,238) /sn:0 /w:[ 0 ]
  //: dip g21 (w11) @(465,123) /sn:0 /w:[ 0 ] /st:1
  //: output g19 (Zero) @(1267,354) /sn:0 /w:[ 1 ]
  mux g32 (.I0(w20), .I1(w11), .S(w15), .Z(w17));   //: @(915,109) /sn:0 /R:1 /w:[ 1 5 1 0 ] /ss:0 /do:0
  not g20 (.I(B), .Z(w12));   //: @(477,207) /sn:0 /w:[ 13 0 ]
  and g15 (.I0(ALU_result), .I1(w1), .Z(Zero));   //: @(1212,354) /sn:0 /w:[ 5 3 0 ]
  add g0 (.A(B), .B(A), .S(w2), .CI(w0), .CO(w4));   //: @(759,286) /sn:0 /R:1 /w:[ 7 5 0 1 0 ]
  //: supply0 g27 (w7) @(651,104) /sn:0 /R:2 /w:[ 1 ]
  tran g13(.Z(w10), .I(ALU_operation[3:0]));   //: @(1016,541) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0

endmodule

module main;    //: root_module
wire [31:0] w4;    //: /sn:0 {0}(388,208)(378,208){1}
wire w3;    //: /sn:0 {0}(388,138)(378,138){1}
wire [31:0] w0;    //: /sn:0 {0}(184,205)(194,205){1}
wire [31:0] w1;    //: /sn:0 {0}(184,139)(194,139){1}
wire [3:0] w2;    //: /sn:0 {0}(279,62)(279,72){1}
//: enddecls

  EXE g0 (.ALU_operation(w2), .A(w1), .B(w0), .ALU_result(w4), .Zero(w3));   //: @(195, 73) /sz:(182, 314) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<1 Ro1<1 ]

endmodule
