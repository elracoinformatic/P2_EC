//: version "1.8.7"

module READ(Read_data_2, Read_register_2, Write_register, mux_RegDst, Read_register_1, Write_data, clk, Sign_ext_32, clr, Sign_ext_in, Read_data_1, RegWrite);
//: interface  /sz:(255, 283) /bd:[ Ti0>RegWrite(135/255) Li0>Sign_ext_in[15:0](237/283) Li1>mux_RegDst(180/283) Li2>Write_register[4:0](151/283) Li3>Read_register_2[4:0](102/283) Li4>Read_register_1[4:0](50/283) Bi0>Write_data[31:0](20/255) Bi1>clr(144/255) Bi2>clk(89/255) Ro0<Sign_ext_out[31:0](250/283) Ro1<Read_data_2[31:0](162/283) Ro2<Read_data_1[31:0](53/283) ]
output [31:0] Read_data_1;    //: /sn:0 /dp:1 {0}(483,82)(616,82)(616,83)(626,83){1}
input [4:0] Write_register;    //: /sn:0 {0}(88,153)(170,153){1}
input [4:0] Read_register_1;    //: /sn:0 /dp:1 {0}(83,67)(334,67){1}
input [4:0] Read_register_2;    //: /sn:0 {0}(334,107)(120,107)(120,131){1}
//: {2}(122,133)(170,133){3}
//: {4}(118,133)(89,133){5}
output [31:0] Read_data_2;    //: /sn:0 /dp:1 {0}(483,174)(561,174)(561,165)(571,165){1}
input [31:0] Write_data;    //: /sn:0 /dp:1 {0}(94,235)(242,235)(242,183)(334,183){1}
input clr;    //: /sn:0 {0}(259,-43)(401,-43)(401,34){1}
input RegWrite;    //: /sn:0 {0}(7,290)(375,290)(375,218){1}
output [31:0] Sign_ext_32;    //: /sn:0 /dp:1 {0}(431,402)(608,402)(608,407)(618,407){1}
input mux_RegDst;    //: /sn:0 {0}(94,210)(186,210)(186,166){1}
input clk;    //: /sn:0 {0}(452,330)(452,264)(443,264)(443,254){1}
input [15:0] Sign_ext_in;    //: /sn:0 {0}(62,401)(316,401)(316,397)(326,397){1}
wire w7;    //: /sn:0 {0}(443,218)(443,238){1}
wire [4:0] w3;    //: /sn:0 /dp:1 {0}(199,143)(334,143){1}
//: enddecls

  BRegs32x32 g4 (.clr(clr), .Read1(Read_register_1), .Read2(Read_register_2), .Write(w3), .WriteData(Write_data), .clk(w7), .RegWrite(RegWrite), .Data1(Read_data_1), .Data2(Read_data_2));   //: @(335, 35) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>0 Li2>1 Li3>1 Bi0>0 Bi1>1 Ro0<0 Ro1<0 ]
  not g8 (.I(clk), .Z(w7));   //: @(443,248) /sn:0 /R:1 /w:[ 1 1 ]
  //: output g16 (Read_data_2) @(568,165) /sn:0 /w:[ 1 ]
  //: input g3 (Read_register_2) @(87,133) /sn:0 /w:[ 5 ]
  //: input g2 (Write_register) @(86,153) /sn:0 /w:[ 0 ]
  //: input g1 (mux_RegDst) @(92,210) /sn:0 /w:[ 0 ]
  signextend g10 (.In(Sign_ext_in), .Out(Sign_ext_32));   //: @(327, 367) /sz:(103, 81) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: input g6 (Read_register_1) @(81,67) /sn:0 /w:[ 0 ]
  //: input g7 (Write_data) @(92,235) /sn:0 /w:[ 0 ]
  //: input g9 (clk) @(452,332) /sn:0 /R:1 /w:[ 0 ]
  //: output g12 (Sign_ext_32) @(615,407) /sn:0 /w:[ 1 ]
  //: input g14 (clr) @(257,-43) /sn:0 /w:[ 0 ]
  //: input g11 (Sign_ext_in) @(60,401) /sn:0 /w:[ 0 ]
  //: joint g5 (Read_register_2) @(120, 133) /w:[ 2 1 4 -1 ]
  //: output g15 (Read_data_1) @(623,83) /sn:0 /w:[ 1 ]
  mux g0 (.I0(Write_register), .I1(Read_register_2), .S(mux_RegDst), .Z(w3));   //: @(186,143) /sn:0 /R:1 /w:[ 1 3 1 0 ] /ss:0 /do:0
  //: input g13 (RegWrite) @(5,290) /sn:0 /w:[ 0 ]

endmodule

module signextend(Out, In);
//: interface  /sz:(183, 170) /bd:[ Li0>In[15:0](65/170) Ro0<Out[31:0](75/170) ]
input [15:0] In;    //: /sn:0 {0}(230,211)(347,211)(347,210)(463,210){1}
//: {2}(464,210)(473,210)(473,302)(614,302){3}
output [31:0] Out;    //: /sn:0 {0}(721,211)(700,211)(700,222)(620,222){1}
wire w3;    //: /sn:0 {0}(614,282)(591,282){1}
//: {2}(587,282)(572,282)(572,264){3}
//: {4}(574,262)(591,262){5}
//: {6}(595,262)(614,262){7}
//: {8}(593,264)(593,272)(614,272){9}
//: {10}(570,262)(538,262)(538,234){11}
//: {12}(540,232)(567,232){13}
//: {14}(571,232)(587,232){15}
//: {16}(591,232)(614,232){17}
//: {18}(589,234)(589,242)(614,242){19}
//: {20}(569,234)(569,252)(614,252){21}
//: {22}(536,232)(529,232)(529,120)(518,120)(518,130){23}
//: {24}(520,132)(532,132){25}
//: {26}(536,132)(542,132)(542,142)(552,142){27}
//: {28}(556,142)(567,142){29}
//: {30}(571,142)(581,142){31}
//: {32}(585,142)(614,142){33}
//: {34}(583,140)(583,130)(598,130)(598,162)(614,162){35}
//: {36}(583,144)(583,152)(614,152){37}
//: {38}(569,144)(569,172)(614,172){39}
//: {40}(554,140)(554,130)(577,130)(577,192)(614,192){41}
//: {42}(554,144)(554,182)(614,182){43}
//: {44}(534,130)(534,120)(549,120)(549,212)(614,212){45}
//: {46}(534,134)(534,202)(614,202){47}
//: {48}(516,132)(464,132)(464,205){49}
//: {50}(518,134)(518,222)(614,222){51}
//: {52}(589,284)(589,292)(614,292){53}
//: enddecls

  //: joint g4 (w3) @(569, 142) /w:[ 30 -1 29 38 ]
  //: joint g8 (w3) @(589, 232) /w:[ 16 -1 15 18 ]
  //: joint g3 (w3) @(583, 142) /w:[ 32 34 31 36 ]
  tran g2(.Z(w3), .I(In[15]));   //: @(464,208) /sn:0 /R:1 /w:[ 49 1 2 ] /ss:0
  concat g1 (.I0(In), .I1(w3), .I2(w3), .I3(w3), .I4(w3), .I5(w3), .I6(w3), .I7(w3), .I8(w3), .I9(w3), .I10(w3), .I11(w3), .I12(w3), .I13(w3), .I14(w3), .I15(w3), .I16(w3), .Z(Out));   //: @(619,222) /sn:0 /w:[ 3 53 0 9 7 21 19 17 51 45 47 41 43 39 35 37 33 1 ] /dr:0
  //: joint g10 (w3) @(538, 232) /w:[ 12 -1 22 11 ]
  //: joint g6 (w3) @(534, 132) /w:[ 26 44 25 46 ]
  //: joint g7 (w3) @(518, 132) /w:[ 24 23 48 50 ]
  //: joint g9 (w3) @(569, 232) /w:[ 14 -1 13 20 ]
  //: joint g12 (w3) @(572, 262) /w:[ 4 -1 10 3 ]
  //: joint g5 (w3) @(554, 142) /w:[ 28 40 27 42 ]
  //: joint g11 (w3) @(593, 262) /w:[ 6 -1 5 8 ]
  //: output g14 (Out) @(718,211) /sn:0 /w:[ 0 ]
  //: input g0 (In) @(228,211) /sn:0 /w:[ 0 ]
  //: joint g13 (w3) @(589, 282) /w:[ 1 -1 2 52 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clk, clr, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>clk(59/69) Li1>RegWr(47/69) Li2>SB[2:0](22/69) Li3>SA[2:0](11/69) Li4>SD[2:0](35/69) Ri0>clr(35/69) Bo0<BOUT[31:0](65/98) Bo1<AOUT[31:0](37/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(207,365)(217,365){1}
wire w7;    //: /sn:0 {0}(353,117)(353,127){1}
wire [31:0] Read_data_1;    //: /sn:0 {0}(484,181)(474,181){1}
wire [4:0] w4;    //: /sn:0 {0}(207,279)(217,279){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(484,290)(474,290){1}
wire [4:0] w3;    //: /sn:0 {0}(207,230)(217,230){1}
wire [31:0] w10;    //: /sn:0 {0}(238,422)(238,412){1}
wire [31:0] w1;    //: /sn:0 {0}(484,378)(474,378){1}
wire w8;    //: /sn:0 {0}(307,422)(307,412){1}
wire [4:0] w2;    //: /sn:0 {0}(207,178)(217,178){1}
wire w5;    //: /sn:0 {0}(207,308)(217,308){1}
wire w9;    //: /sn:0 {0}(362,422)(362,412){1}
//: enddecls

  READ g0 (.RegWrite(w7), .Sign_ext_in(w6), .mux_RegDst(w5), .Write_register(w4), .Read_register_2(w3), .Read_register_1(w2), .Write_data(w10), .clr(w9), .clk(w8), .Sign_ext_out(w1), .Read_data_2(w0), .Read_data_1(Read_data_1));   //: @(218, 128) /sz:(255, 283) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Bi0>1 Bi1>1 Bi2>1 Ro0<1 Ro1<1 Ro2<1 ]

endmodule
