//: version "1.8.7"

module MEM(write_data, MemRead, memWrite, read_data, Address);
//: interface  /sz:(128, 174) /bd:[ Ti0>memWrite(62/128) Li0>Address[31:0](43/174) Li1>write_data[31:0](112/174) Bi0>MemRead(59/128) Ro0<read_data[31:0](35/174) ]
input [31:0] write_data;    //: /sn:0 {0}(316,166)(458,166)(458,192)(488,192){1}
output [31:0] read_data;    //: /sn:0 /dp:1 {0}(504,192)(514,192)(514,247){1}
//: {2}(516,249)(545,249){3}
//: {4}(512,249)(443,249){5}
input memWrite;    //: /sn:0 {0}(317,198)(329,198){1}
//: {2}(333,198)(379,198){3}
//: {4}(383,198)(392,198){5}
//: {6}(381,196)(381,111)(496,111)(496,187){7}
//: {8}(331,200)(331,228)(312,228)(312,244)(282,244)(282,307)(311,307){9}
input MemRead;    //: /sn:0 {0}(304,386)(329,386)(329,384){1}
//: {2}(331,382)(341,382)(341,386)(375,386){3}
//: {4}(329,380)(329,325)(301,325)(301,312)(311,312){5}
input [31:0] Address;    //: /sn:0 {0}(379,251)(408,251){1}
wire w4;    //: /sn:0 {0}(408,198)(426,198)(426,226){1}
wire w3;    //: /sn:0 {0}(391,386)(433,386)(433,276){1}
wire w2;    //: /sn:0 {0}(332,310)(419,310)(419,276){1}
//: enddecls

  //: input g8 (write_data) @(314,166) /sn:0 /w:[ 0 ]
  //: input g4 (MemRead) @(302,386) /sn:0 /w:[ 0 ]
  //: input g3 (memWrite) @(315,198) /sn:0 /w:[ 0 ]
  //: output g2 (read_data) @(542,249) /sn:0 /w:[ 3 ]
  //: input g1 (Address) @(377,251) /sn:0 /w:[ 0 ]
  not g10 (.I(MemRead), .Z(w3));   //: @(381,386) /sn:0 /w:[ 3 0 ]
  //: joint g6 (read_data) @(514, 249) /w:[ 2 1 4 -1 ]
  not g7 (.I(memWrite), .Z(w4));   //: @(398,198) /sn:0 /w:[ 5 0 ]
  nor g9 (.I0(memWrite), .I1(MemRead), .Z(w2));   //: @(322,310) /sn:0 /w:[ 9 5 0 ]
  //: joint g12 (MemRead) @(329, 382) /w:[ 2 4 -1 1 ]
  //: joint g11 (memWrite) @(331, 198) /w:[ 2 -1 1 8 ]
  bufif1 g5 (.Z(read_data), .I(write_data), .E(memWrite));   //: @(494,192) /sn:0 /w:[ 0 1 7 ]
  ram g0 (.A(Address), .D(read_data), .WE(w4), .OE(w3), .CS(w2));   //: @(426,250) /sn:0 /w:[ 1 5 1 1 1 ]
  //: joint g13 (memWrite) @(381, 198) /w:[ 4 6 3 -1 ]

endmodule

module ALUCtrl(ALUOp, ALUCtrl, funct);
//: interface  /sz:(171, 213) /bd:[ Li0>ALUOp[1:0](35/213) Li1>funct[5:0](103/213) Ro0<ALUCtrl[3:0](50/213) ]
output [3:0] ALUCtrl;    //: /sn:0 /dp:1 {0}(1002,416)(1057,416)(1057,423)(1106,423){1}
supply0 [3:0] w4;    //: /sn:0 {0}(839,369)(839,398)(973,398){1}
supply0 w3;    //: /sn:0 {0}(610,456)(610,454)(611,454)(611,444){1}
input [1:0] ALUOp;    //: /sn:0 {0}(314,545)(989,545)(989,439){1}
input [5:0] funct;    //: /sn:0 {0}(407,426)(527,426)(527,419)(593,419){1}
wire [3:0] w0;    //: /sn:0 {0}(723,451)(881,451)(881,422)(973,422){1}
wire [3:0] w1;    //: /sn:0 {0}(628,417)(804,417)(804,410)(973,410){1}
wire [3:0] w2;    //: /sn:0 {0}(822,482)(963,482)(963,434)(973,434){1}
//: enddecls

  //: input g4 (ALUOp) @(312,545) /sn:0 /w:[ 0 ]
  //: output g8 (ALUCtrl) @(1103,423) /sn:0 /w:[ 1 ]
  mux g3 (.I0(w2), .I1(w0), .I2(w1), .I3(w4), .S(ALUOp), .Z(ALUCtrl));   //: @(989,416) /sn:0 /R:1 /w:[ 1 1 1 1 1 0 ] /ss:0 /do:0
  //: input g2 (funct) @(405,426) /sn:0 /w:[ 0 ]
  //: supply0 g1 (w3) @(610,462) /sn:0 /w:[ 0 ]
  //: dip g6 (w0) @(685,451) /sn:0 /R:1 /w:[ 0 ] /st:6
  //: supply0 g7 (w4) @(839,363) /sn:0 /R:2 /w:[ 0 ]
  //: dip g5 (w2) @(784,482) /sn:0 /R:1 /w:[ 0 ] /st:2
  rom g0 (.A(funct), .D(w1), .OE(w3));   //: @(611,418) /sn:0 /w:[ 1 0 1 ]

endmodule

module ctrl(RegDst, ALUSrc, instruction, MemRead, Jump, MemtoReg, Branch, RegWrite, MemWrite, ALUOp);
//: interface  /sz:(171, 276) /bd:[ Li0>instruction[5:0](47/276) Ro0<RegWrite(240/276) Ro1<ALUSrc(211/276) Ro2<MemWrite(175/276) Ro3<MemtoReg(120/276) Ro4<ALUOp[1:0](151/276) Ro5<MemRead(91/276) Ro6<Branch(67/276) Ro7<Jump(42/276) Ro8<RegDst(22/276) ]
output Branch;    //: /sn:0 {0}(432,-28)(561,-28){1}
supply0 w3;    //: /sn:0 {0}(309,8)(309,-50)(331,-50)(331,-60){1}
output MemWrite;    //: /sn:0 {0}(432,193)(440,193)(440,194)(565,194){1}
output ALUSrc;    //: /sn:0 {0}(432,227)(440,227)(440,228)(588,228){1}
input [5:0] instruction;    //: /sn:0 {0}(21,-73)(303,-73)(303,-85)(313,-85){1}
output RegDst;    //: /sn:0 {0}(432,-62)(558,-62){1}
output RegWrite;    //: /sn:0 {0}(432,259)(440,259)(440,258)(585,258){1}
output [1:0] ALUOp;    //: /sn:0 {0}(432,144)(440,144)(440,145)(577,145){1}
output MemtoReg;    //: /sn:0 {0}(433,86)(441,86)(441,94)(563,94){1}
output MemRead;    //: /sn:0 {0}(432,43)(440,43)(440,48)(566,48){1}
output Jump;    //: /sn:0 {0}(432,9)(440,9)(440,12)(563,12){1}
wire [9:0] w1;    //: /sn:0 {0}(348,-87)(428,-87)(428,-63){1}
//: {2}(428,-62)(428,-29){3}
//: {4}(428,-28)(428,8){5}
//: {6}(428,9)(428,42){7}
//: {8}(428,43)(428,63)(429,63)(429,85){9}
//: {10}(429,86)(429,133)(428,133)(428,143){11}
//: {12}(428,144)(428,192){13}
//: {14}(428,193)(428,226){15}
//: {16}(428,227)(428,258){17}
//: {18}(428,259)(428,412){19}
//: enddecls

  tran g8(.Z(Jump), .I(w1[7]));   //: @(426,9) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  tran g4(.Z(RegDst), .I(w1[9]));   //: @(426,-62) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: output g3 (RegDst) @(555,-62) /sn:0 /w:[ 1 ]
  tran g16(.Z(MemWrite), .I(w1[2]));   //: @(426,193) /sn:0 /R:2 /w:[ 0 14 13 ] /ss:1
  //: output g17 (ALUSrc) @(585,228) /sn:0 /w:[ 1 ]
  //: input g2 (instruction) @(19,-73) /sn:0 /w:[ 0 ]
  //: supply0 g1 (w3) @(309,14) /sn:0 /w:[ 0 ]
  tran g18(.Z(ALUSrc), .I(w1[1]));   //: @(426,227) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  tran g10(.Z(MemRead), .I(w1[6]));   //: @(426,43) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  tran g6(.Z(Branch), .I(w1[8]));   //: @(426,-28) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: output g9 (MemRead) @(563,48) /sn:0 /w:[ 1 ]
  //: output g7 (Jump) @(560,12) /sn:0 /w:[ 1 ]
  tran g12(.Z(MemtoReg), .I(w1[5]));   //: @(427,86) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  //: output g11 (MemtoReg) @(560,94) /sn:0 /w:[ 1 ]
  //: output g5 (Branch) @(558,-28) /sn:0 /w:[ 1 ]
  tran g14(.Z(ALUOp), .I(w1[4:3]));   //: @(426,144) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  //: output g19 (RegWrite) @(582,258) /sn:0 /w:[ 1 ]
  tran g20(.Z(RegWrite), .I(w1[0]));   //: @(426,259) /sn:0 /R:2 /w:[ 0 18 17 ] /ss:1
  rom g0 (.A(instruction), .D(w1), .OE(w3));   //: @(331,-86) /sn:0 /w:[ 1 0 1 ]
  //: output g15 (MemWrite) @(562,194) /sn:0 /w:[ 1 ]
  //: output g13 (ALUOp) @(574,145) /sn:0 /w:[ 1 ]

endmodule

module READ(Read_register_2, Read_data_2, Write_register, mux_RegDst, Read_register_1, clk, Write_data, Sign_ext_out, Sign_ext_in, clr, Read_data_1, RegWrite);
//: interface  /sz:(255, 283) /bd:[ Ti0>RegWrite(135/255) Li0>Read_register_1[4:0](50/283) Li1>Read_register_2[4:0](102/283) Li2>Write_register[4:0](151/283) Li3>mux_RegDst(180/283) Li4>Sign_ext_in[15:0](237/283) Bi0>clk(89/255) Bi1>clr(144/255) Bi2>Write_data[31:0](20/255) Ro0<Read_data_1[31:0](53/283) Ro1<Read_data_2[31:0](162/283) Ro2<Sign_ext_out[31:0](250/283) ]
output [31:0] Read_data_1;    //: /sn:0 /dp:1 {0}(483,82)(616,82)(616,83)(626,83){1}
input [4:0] Write_register;    //: /sn:0 {0}(66,173)(150,173)(150,133)(170,133){1}
input [4:0] Read_register_1;    //: /sn:0 /dp:1 {0}(83,67)(334,67){1}
input [4:0] Read_register_2;    //: /sn:0 /dp:1 {0}(89,133)(118,133){1}
//: {2}(120,131)(120,107)(334,107){3}
//: {4}(120,135)(120,153)(170,153){5}
output [31:0] Read_data_2;    //: /sn:0 /dp:1 {0}(483,174)(561,174)(561,165)(571,165){1}
input [31:0] Write_data;    //: /sn:0 /dp:1 {0}(94,235)(242,235)(242,183)(334,183){1}
input RegWrite;    //: /sn:0 {0}(7,290)(375,290)(375,218){1}
input clr;    //: /sn:0 {0}(259,-43)(401,-43)(401,34){1}
input mux_RegDst;    //: /sn:0 {0}(94,210)(186,210)(186,166){1}
input clk;    //: /sn:0 {0}(452,330)(452,264)(443,264)(443,254){1}
output [31:0] Sign_ext_out;    //: /sn:0 /dp:1 {0}(420,408)(597,408)(597,407)(618,407){1}
input [15:0] Sign_ext_in;    //: /sn:0 {0}(62,401)(305,401)(305,403)(315,403){1}
wire w7;    //: /sn:0 {0}(443,218)(443,238){1}
wire [4:0] w3;    //: /sn:0 /dp:1 {0}(199,143)(334,143){1}
//: enddecls

  not g8 (.I(clk), .Z(w7));   //: @(443,248) /sn:0 /R:1 /w:[ 1 1 ]
  BRegs32x32 g4 (.clr(clr), .Read1(Read_register_1), .Read2(Read_register_2), .Write(w3), .WriteData(Write_data), .clk(w7), .RegWrite(RegWrite), .Data1(Read_data_1), .Data2(Read_data_2));   //: @(335, 35) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>1 Li3>1 Bi0>0 Bi1>1 Ro0<0 Ro1<0 ]
  //: input g3 (Read_register_2) @(87,133) /sn:0 /w:[ 0 ]
  //: output g16 (Read_data_2) @(568,165) /sn:0 /w:[ 1 ]
  //: input g2 (Write_register) @(64,173) /sn:0 /w:[ 0 ]
  //: input g1 (mux_RegDst) @(92,210) /sn:0 /w:[ 0 ]
  signextend g10 (.In(Sign_ext_in), .Out(Sign_ext_out));   //: @(316, 373) /sz:(103, 81) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: input g6 (Read_register_1) @(81,67) /sn:0 /w:[ 0 ]
  //: input g9 (clk) @(452,332) /sn:0 /R:1 /w:[ 0 ]
  //: input g7 (Write_data) @(92,235) /sn:0 /w:[ 0 ]
  //: output g12 (Sign_ext_out) @(615,407) /sn:0 /w:[ 1 ]
  //: joint g5 (Read_register_2) @(120, 133) /w:[ -1 2 1 4 ]
  //: input g11 (Sign_ext_in) @(60,401) /sn:0 /w:[ 0 ]
  //: input g14 (clr) @(257,-43) /sn:0 /w:[ 0 ]
  mux g0 (.I0(Read_register_2), .I1(Write_register), .S(mux_RegDst), .Z(w3));   //: @(186,143) /sn:0 /R:1 /w:[ 5 1 1 0 ] /ss:0 /do:0
  //: output g15 (Read_data_1) @(623,83) /sn:0 /w:[ 1 ]
  //: input g13 (RegWrite) @(5,290) /sn:0 /w:[ 0 ]

endmodule

module signextend(Out, In);
//: interface  /sz:(183, 170) /bd:[ Li0>In[15:0](65/170) Ro0<Out[31:0](75/170) ]
input [15:0] In;    //: /sn:0 {0}(230,211)(347,211)(347,210)(463,210){1}
//: {2}(464,210)(473,210)(473,302)(614,302){3}
output [31:0] Out;    //: /sn:0 {0}(721,211)(700,211)(700,222)(620,222){1}
wire w3;    //: /sn:0 {0}(614,282)(591,282){1}
//: {2}(587,282)(572,282)(572,264){3}
//: {4}(574,262)(591,262){5}
//: {6}(595,262)(614,262){7}
//: {8}(593,264)(593,272)(614,272){9}
//: {10}(570,262)(538,262)(538,234){11}
//: {12}(540,232)(567,232){13}
//: {14}(571,232)(587,232){15}
//: {16}(591,232)(614,232){17}
//: {18}(589,234)(589,242)(614,242){19}
//: {20}(569,234)(569,252)(614,252){21}
//: {22}(536,232)(529,232)(529,120)(518,120)(518,130){23}
//: {24}(520,132)(532,132){25}
//: {26}(536,132)(542,132)(542,142)(552,142){27}
//: {28}(556,142)(567,142){29}
//: {30}(571,142)(581,142){31}
//: {32}(585,142)(614,142){33}
//: {34}(583,140)(583,130)(598,130)(598,162)(614,162){35}
//: {36}(583,144)(583,152)(614,152){37}
//: {38}(569,144)(569,172)(614,172){39}
//: {40}(554,140)(554,130)(577,130)(577,192)(614,192){41}
//: {42}(554,144)(554,182)(614,182){43}
//: {44}(534,130)(534,120)(549,120)(549,212)(614,212){45}
//: {46}(534,134)(534,202)(614,202){47}
//: {48}(516,132)(464,132)(464,205){49}
//: {50}(518,134)(518,222)(614,222){51}
//: {52}(589,284)(589,292)(614,292){53}
//: enddecls

  //: joint g8 (w3) @(589, 232) /w:[ 16 -1 15 18 ]
  //: joint g4 (w3) @(569, 142) /w:[ 30 -1 29 38 ]
  //: joint g3 (w3) @(583, 142) /w:[ 32 34 31 36 ]
  tran g2(.Z(w3), .I(In[15]));   //: @(464,208) /sn:0 /R:1 /w:[ 49 1 2 ] /ss:0
  concat g1 (.I0(In), .I1(w3), .I2(w3), .I3(w3), .I4(w3), .I5(w3), .I6(w3), .I7(w3), .I8(w3), .I9(w3), .I10(w3), .I11(w3), .I12(w3), .I13(w3), .I14(w3), .I15(w3), .I16(w3), .Z(Out));   //: @(619,222) /sn:0 /w:[ 3 53 0 9 7 21 19 17 51 45 47 41 43 39 35 37 33 1 ] /dr:0
  //: joint g10 (w3) @(538, 232) /w:[ 12 -1 22 11 ]
  //: joint g6 (w3) @(534, 132) /w:[ 26 44 25 46 ]
  //: joint g9 (w3) @(569, 232) /w:[ 14 -1 13 20 ]
  //: joint g7 (w3) @(518, 132) /w:[ 24 23 48 50 ]
  //: joint g12 (w3) @(572, 262) /w:[ 4 -1 10 3 ]
  //: output g14 (Out) @(718,211) /sn:0 /w:[ 0 ]
  //: joint g11 (w3) @(593, 262) /w:[ 6 -1 5 8 ]
  //: joint g5 (w3) @(554, 142) /w:[ 28 40 27 42 ]
  //: input g0 (In) @(228,211) /sn:0 /w:[ 0 ]
  //: joint g13 (w3) @(589, 282) /w:[ 1 -1 2 52 ]

endmodule

module fetch(reset, clk, Inst, PCNext, PCNew);
//: interface  /sz:(420, 354) /bd:[ Li0>PCNew[31:0](181/354) Li1>reset(96/354) Li2>clk(262/354) Ro0<Inst[31:0](271/354) Ro1<PCNext[31:0](49/354) ]
supply0 w4;    //: /sn:0 {0}(258,62)(258,93)(257,93)(257,101){1}
input [31:0] PCNew;    //: /sn:0 {0}(241,139)(231,139)(231,138)(163,138){1}
output [31:0] Inst;    //: /sn:0 /dp:1 {0}(366,149)(468,149)(468,137)(574,137){1}
output [31:0] PCNext;    //: /sn:0 /dp:1 {0}(436,68)(541,68)(541,65)(551,65){1}
supply0 w1;    //: /sn:0 {0}(353,202)(353,195)(349,195)(349,176){1}
input clk;    //: /sn:0 {0}(139,189)(252,189)(252,177){1}
supply0 w2;    //: /sn:0 {0}(419,-6)(419,37)(421,37)(421,44){1}
input reset;    //: /sn:0 {0}(151,75)(247,75)(247,101){1}
wire w7;    //: /sn:0 {0}(421,92)(421,121){1}
wire [31:0] w0;    //: /sn:0 {0}(262,139)(289,139){1}
//: {2}(293,139)(310,139)(310,151)(331,151){3}
//: {4}(291,137)(291,52)(407,52){5}
wire [31:0] w3;    //: /sn:0 {0}(382,80)(397,80)(397,84)(407,84){1}
//: enddecls

  add g8 (.A(w3), .B(w0), .S(PCNext), .CI(w2), .CO(w7));   //: @(423,68) /sn:0 /R:1 /w:[ 1 5 0 1 0 ]
  rom Imemo (.A(w0), .D(Inst), .OE(w1));   //: @(349,150) /w:[ 3 0 1 ]
  register g3 (.Q(w0), .D(PCNew), .EN(w4), .CLR(reset), .CK(clk));   //: @(252,139) /sn:0 /R:1 /w:[ 0 0 1 1 1 ]
  //: input g2 (reset) @(149,75) /sn:0 /w:[ 0 ]
  //: input g1 (clk) @(137,189) /sn:0 /w:[ 0 ]
  //: dip g10 (w3) @(344,80) /sn:0 /R:1 /w:[ 0 ] /st:1
  //: output g6 (Inst) @(571,137) /sn:0 /w:[ 1 ]
  //: supply0 g7 (w4) @(258,56) /sn:0 /R:2 /w:[ 0 ]
  //: joint g9 (w0) @(291, 139) /w:[ 2 4 1 -1 ]
  //: supply0 g12 (w2) @(419,-12) /sn:0 /R:2 /w:[ 0 ]
  //: supply0 g5 (w1) @(353,208) /sn:0 /w:[ 0 ]
  //: output g11 (PCNext) @(548,65) /sn:0 /w:[ 1 ]
  //: input g0 (PCNew) @(161,138) /sn:0 /w:[ 1 ]

endmodule

module ALU(Zero_signal, B, ALU_operation, A, ALU_result);
//: interface  /sz:(127, 166) /bd:[ Ti0>ALU_operation[3:0](64/127) Li0>A[31:0](46/166) Li1>B[31:0](108/166) Ro0<Zero(52/166) Ro1<ALU_result[31:0](106/166) ]
input [31:0] B;    //: /sn:0 {0}(415,270)(468,270){1}
//: {2}(472,270)(594,270){3}
//: {4}(598,270)(643,270){5}
//: {6}(647,270)(700,270)(700,302)(743,302){7}
//: {8}(645,272)(645,370)(720,370){9}
//: {10}(596,272)(596,392)(718,392){11}
//: {12}(470,268)(470,207)(471,207){13}
supply0 w7;    //: /sn:0 /dp:1 {0}(651,129)(651,110){1}
output [31:0] ALU_result;    //: /sn:0 /dp:1 {0}(1029,324)(1108,324){1}
//: {2}(1112,324)(1147,324)(1147,292)(1194,292){3}
//: {4}(1110,326)(1110,363)(1134,363){5}
input [31:0] A;    //: /sn:0 {0}(412,238)(610,238){1}
//: {2}(614,238)(659,238){3}
//: {4}(663,238)(708,238)(708,270)(743,270){5}
//: {6}(661,240)(661,365)(720,365){7}
//: {8}(612,236)(612,137)(637,137){9}
//: {10}(612,240)(612,387)(718,387){11}
supply0 w0;    //: /sn:0 {0}(757,243)(757,262){1}
supply0 w3;    //: /sn:0 /dp:1 {0}(552,145)(552,123){1}
supply0 [31:0] w20;    //: /sn:0 {0}(805,115)(805,119)(899,119){1}
input [3:0] ALU_operation;    //: /sn:0 {0}(428,544)(723,544)(723,543)(1016,543){1}
//: {2}(1017,543)(1078,543){3}
output Zero_signal;    //: /sn:0 /dp:1 {0}(1219,391)(1342,391)(1342,388)(1352,388){1}
supply0 [31:0] w5;    //: /sn:0 {0}(825,318)(857,318)(857,317)(867,317){1}
//: {2}(869,315)(869,314)(1000,314){3}
//: {4}(869,319)(869,320)(983,320){5}
//: {6}(987,320)(1000,320){7}
//: {8}(985,322)(985,327)(1000,327){9}
wire [31:0] w6;    //: /sn:0 {0}(567,169)(637,169){1}
wire [31:0] w16;    //: /sn:0 {0}(666,153)(818,153)(818,159){1}
//: {2}(818,160)(818,307)(1000,307){3}
wire Zero;    //: /sn:0 /dp:1 {0}(822,160)(915,160)(915,132){1}
wire w4;    //: /sn:0 {0}(757,310)(757,338){1}
wire [31:0] w18;    //: /sn:0 {0}(741,368)(793,368)(793,347)(1000,347){1}
wire [31:0] w12;    //: /sn:0 {0}(487,207)(512,207)(512,185)(538,185){1}
wire w19;    //: /sn:0 {0}(651,177)(651,197){1}
wire [2:0] w10;    //: /sn:0 {0}(1017,538)(1017,442)(1016,442)(1016,347){1}
wire w8;    //: /sn:0 {0}(552,193)(552,203)(565,203)(565,213){1}
wire [31:0] w17;    //: /sn:0 {0}(928,109)(990,109)(990,300)(1000,300){1}
wire w14;    //: /sn:0 {0}(1155,363)(1193,363)(1193,391)(1203,391){1}
wire [31:0] w2;    //: /sn:0 {0}(772,286)(800,286)(800,334)(1000,334){1}
wire [31:0] w11;    //: /sn:0 {0}(465,133)(465,153)(518,153){1}
//: {2}(522,153)(538,153){3}
//: {4}(520,151)(520,99)(899,99){5}
wire [31:0] w9;    //: /sn:0 {0}(739,390)(803,390)(803,340)(1000,340){1}
//: enddecls

  or g4 (.I0(A), .I1(B), .Z(w9));   //: @(729,390) /sn:0 /w:[ 11 11 0 ]
  //: joint g8 (A) @(612, 238) /w:[ 2 8 1 10 ]
  and g3 (.I0(A), .I1(B), .Z(w18));   //: @(731,368) /sn:0 /w:[ 7 9 0 ]
  //: supply0 g16 (w5) @(819,318) /sn:0 /R:3 /w:[ 0 ]
  not g17 (.I(w14), .Z(Zero_signal));   //: @(1209,391) /sn:0 /w:[ 1 0 ]
  add g26 (.A(w6), .B(A), .S(w16), .CI(w7), .CO(w19));   //: @(653,153) /sn:0 /R:1 /w:[ 1 9 0 0 0 ]
  or g2 (.I0(ALU_result), .Z(w14));   //: @(1145,363) /sn:0 /w:[ 5 0 ]
  //: joint g23 (B) @(470, 270) /w:[ 2 12 1 -1 ]
  //: joint g30 (w5) @(869, 317) /w:[ -1 2 1 4 ]
  //: joint g1 (A) @(661, 238) /w:[ 4 -1 3 6 ]
  //: supply0 g24 (w3) @(552,117) /sn:0 /R:2 /w:[ 1 ]
  mux g29 (.I0(w18), .I1(w9), .I2(w2), .I3(w5), .I4(w5), .I5(w5), .I6(w16), .I7(w17), .S(w10), .Z(ALU_result));   //: @(1016,324) /sn:0 /R:1 /w:[ 1 1 1 9 7 3 3 1 1 0 ] /ss:0 /do:0
  //: output g18 (Zero_signal) @(1349,388) /sn:0 /w:[ 1 ]
  //: supply0 g10 (w0) @(757,237) /sn:0 /R:2 /w:[ 0 ]
  led g25 (.I(w8));   //: @(565,220) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: input g6 (B) @(413,270) /sn:0 /w:[ 0 ]
  //: joint g7 (B) @(645, 270) /w:[ 6 -1 5 8 ]
  //: joint g9 (B) @(596, 270) /w:[ 4 -1 3 10 ]
  //: joint g35 (w11) @(520, 153) /w:[ 2 4 1 -1 ]
  add g22 (.A(w12), .B(w11), .S(w6), .CI(w3), .CO(w8));   //: @(554,169) /sn:0 /R:1 /w:[ 1 3 0 0 0 ]
  //: joint g31 (w5) @(985, 320) /w:[ 6 -1 5 8 ]
  tran g33(.Z(Zero), .I(w16[31]));   //: @(816,160) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: input g12 (ALU_operation) @(426,544) /sn:0 /w:[ 0 ]
  led g28 (.I(w19));   //: @(651,204) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: supply0 g34 (w20) @(805,109) /sn:0 /R:2 /w:[ 0 ]
  //: input g5 (A) @(410,238) /sn:0 /w:[ 0 ]
  led g11 (.I(w4));   //: @(757,345) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: output g14 (ALU_result) @(1191,292) /sn:0 /w:[ 3 ]
  //: dip g21 (w11) @(465,123) /sn:0 /w:[ 0 ] /st:1
  not g20 (.I(B), .Z(w12));   //: @(477,207) /sn:0 /w:[ 13 0 ]
  mux g32 (.I0(w20), .I1(w11), .S(Zero), .Z(w17));   //: @(915,109) /sn:0 /R:1 /w:[ 1 5 1 0 ] /ss:0 /do:0
  //: joint g15 (ALU_result) @(1110, 324) /w:[ 2 -1 1 4 ]
  add g0 (.A(B), .B(A), .S(w2), .CI(w0), .CO(w4));   //: @(759,286) /sn:0 /R:1 /w:[ 7 5 0 1 0 ]
  //: supply0 g27 (w7) @(651,104) /sn:0 /R:2 /w:[ 1 ]
  tran g13(.Z(w10), .I(ALU_operation[2:0]));   //: @(1017,541) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0

endmodule

module EXE(ALU_result, Zero_signal, data_read_2, data_read_1, INM32, PCNext, branch_target, ALU_operation);
//: interface  /sz:(185, 314) /bd:[ Ti0>ALU_operation[3:0](85/185) Li0>data_read_2[31:0](272/314) Li1>data_read_1[31:0](239/314) Li2>PCNext[31:0](91/314) Li3>INM32[31:0](126/314) Ro0<Zero_signal(242/314) Ro1<ALU_result[31:0](283/314) Ro2<branch_target[31:0](90/314) ]
output [31:0] ALU_result;    //: /sn:0 {0}(540,374)(679,374){1}
input [3:0] ALU_operation;    //: /sn:0 {0}(406,120)(464,120)(464,244){1}
input [31:0] data_read_2;    //: /sn:0 {0}(166,377)(387,377){1}
input [31:0] PCNext;    //: /sn:0 {0}(113,514)(431,514)(431,571)(441,571){1}
output Zero_signal;    //: /sn:0 {0}(540,308)(675,308){1}
output [31:0] branch_target;    //: /sn:0 /dp:1 {0}(470,587)(550,587)(550,586)(560,586){1}
input [31:0] INM32;    //: /sn:0 /dp:1 {0}(116,623)(431,623)(431,603)(441,603){1}
supply0 w5;    //: /sn:0 {0}(455,524)(455,563){1}
input [31:0] data_read_1;    //: /sn:0 {0}(170,301)(387,301){1}
wire w3;    //: /sn:0 /dp:1 {0}(455,647)(455,611){1}
//: enddecls

  led g8 (.I(w3));   //: @(455,654) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: output g4 (ALU_result) @(676,374) /sn:0 /w:[ 1 ]
  //: output g3 (Zero_signal) @(672,308) /sn:0 /w:[ 1 ]
  //: input g2 (data_read_2) @(164,377) /sn:0 /w:[ 0 ]
  //: input g1 (data_read_1) @(168,301) /sn:0 /w:[ 0 ]
  //: input g10 (INM32) @(114,623) /sn:0 /w:[ 0 ]
  add g6 (.A(INM32), .B(PCNext), .S(branch_target), .CI(w5), .CO(w3));   //: @(457,587) /sn:0 /R:1 /w:[ 1 1 0 1 1 ]
  //: input g9 (PCNext) @(111,514) /sn:0 /w:[ 0 ]
  //: supply0 g7 (w5) @(455,518) /sn:0 /R:2 /w:[ 0 ]
  //: output g11 (branch_target) @(557,586) /sn:0 /w:[ 1 ]
  //: input g5 (ALU_operation) @(404,120) /sn:0 /w:[ 0 ]
  ALU g0 (.ALU_operation(ALU_operation), .B(data_read_2), .A(data_read_1), .ALU_result(ALU_result), .Zero_signal(Zero_signal));   //: @(388, 245) /sz:(151, 203) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<0 Ro1<0 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Li0>WriteData[31:0](148/182) Li1>Write[4:0](108/182) Li2>Read2[4:0](72/182) Li3>Read1[4:0](32/182) Bi0>RegWrite(40/147) Bi1>clk(108/147) Ro0<Data2[31:0](139/182) Ro1<Data1[31:0](47/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clr, clk, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>SD[2:0](35/69) Li1>SA[2:0](11/69) Li2>SB[2:0](22/69) Li3>RegWr(47/69) Li4>clk(59/69) Ri0>clr(35/69) Bo0<AOUT[31:0](37/98) Bo1<BOUT[31:0](65/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(403,572)(316,572)(316,571)(307,571){1}
wire w13;    //: /sn:0 {0}(491,619)(491,669)(-146,669)(-146,465){1}
//: {2}(-144,463)(-71,463)(-71,453)(-63,453){3}
//: {4}(-148,463)(-240,463){5}
wire [31:0] w16;    //: /sn:0 {0}(660,388)(828,388)(828,325)(866,325){1}
wire [31:0] w4;    //: /sn:0 {0}(78,468)(86,468)(86,429)(183,429){1}
//: {2}(184,429)(207,429)(207,431)(231,431){3}
//: {4}(232,431)(242,431)(242,446)(190,446)(190,496)(146,496)(146,484)(143,484){5}
//: {6}(142,484)(116,484)(116,520)(249,520){7}
//: {8}(250,520)(259,520)(259,514)(295,514){9}
//: {10}(296,514)(331,514)(331,507)(343,507){11}
//: {12}(344,507)(354,507)(354,516)(343,516)(343,528)(321,528)(321,546)(303,546)(303,570){13}
//: {14}(303,571)(303,627){15}
wire [31:0] w25;    //: /sn:0 /dp:1 {0}(817,433)(719,433){1}
//: {2}(717,431)(717,421)(737,421)(737,212)(866,212){3}
//: {4}(717,435)(717,585)(660,585){5}
wire w39;    //: /sn:0 {0}(428,-2)(1323,-2)(1323,252)(1378,252)(1378,242){1}
wire [31:0] w3;    //: /sn:0 {0}(78,261)(130,261)(130,189)(545,189){1}
//: {2}(546,189)(827,189)(827,179){3}
//: {4}(829,177)(866,177){5}
//: {6}(827,175)(827,-32)(1106,-32){7}
wire [31:0] w22;    //: /sn:0 {0}(1053,176)(1096,176)(1096,-52)(1106,-52){1}
wire w36;    //: /sn:0 {0}(428,-41)(999,-41)(999,56)(1065,56){1}
wire w0;    //: /sn:0 {0}(-232,690)(548,690)(548,619){1}
wire [27:0] w29;    //: /sn:0 {0}(232,426)(232,155)(628,155){1}
wire [31:0] w30;    //: /sn:0 {0}(634,160)(683,160)(683,-81)(1154,-81)(1154,-72)(1194,-72){1}
wire w37;    //: /sn:0 {0}(428,-23)(1443,-23)(1443,322)(1224,322)(1224,312){1}
wire w42;    //: /sn:0 {0}(428,87)(539,87)(539,334){1}
wire [3:0] w19;    //: /sn:0 {0}(546,184)(546,165)(628,165){1}
wire w18;    //: /sn:0 {0}(1086,59)(1122,59)(1122,-19){1}
wire [4:0] w10;    //: /sn:0 {0}(403,385)(250,385)(250,515){1}
wire [31:0] w23;    //: /sn:0 {0}(1053,369)(1116,369)(1116,234){1}
//: {2}(1118,232)(1141,232)(1141,340)(1311,340)(1311,229)(1362,229){3}
//: {4}(1116,230)(1116,180)(1164,180){5}
wire w24;    //: /sn:0 {0}(1053,328)(1061,328)(1061,61)(1065,61){1}
wire w1;    //: /sn:0 {0}(-63,303)(-73,303){1}
wire [31:0] w31;    //: /sn:0 {0}(846,443)(856,443)(856,358)(866,358){1}
wire [31:0] w32;    //: /sn:0 {0}(1391,219)(1401,219)(1401,644)(424,644)(424,619){1}
wire [4:0] w8;    //: /sn:0 {0}(403,486)(344,486)(344,502){1}
wire [1:0] w44;    //: /sn:0 {0}(680,-250)(629,-250)(629,21)(428,21){1}
wire [31:0] w33;    //: /sn:0 {0}(1135,-42)(1184,-42)(1184,-52)(1194,-52){1}
wire [31:0] w28;    //: /sn:0 {0}(1294,164)(1352,164)(1352,209)(1362,209){1}
wire [31:0] w35;    //: /sn:0 {0}(1223,-62)(1239,-62)(1239,-155)(-73,-155)(-73,380)(-63,380){1}
wire w14;    //: /sn:0 {0}(428,-59)(1081,-59)(1081,-136)(1179,-136)(1179,-29)(1210,-29)(1210,-39){1}
wire [3:0] w45;    //: /sn:0 {0}(816,-243)(952,-243)(952,85){1}
wire [5:0] w2;    //: /sn:0 {0}(255,-56)(143,-56)(143,479){1}
wire w11;    //: /sn:0 {0}(428,-74)(456,-74)(456,306)(381,306)(381,515)(403,515){1}
wire w41;    //: /sn:0 {0}(428,65)(800,65)(800,476)(833,476)(833,466){1}
wire [31:0] w15;    //: /sn:0 {0}(660,497)(785,497){1}
//: {2}(789,497)(1156,497)(1156,249)(1164,249){3}
//: {4}(787,495)(787,453)(817,453){5}
wire [5:0] w43;    //: /sn:0 {0}(680,-216)(184,-216)(184,424){1}
wire [4:0] w9;    //: /sn:0 {0}(403,437)(296,437)(296,509){1}
wire w40;    //: /sn:0 {0}(428,39)(1227,39)(1227,136){1}
//: enddecls

  concat g4 (.I0(w19), .I1(w29), .Z(w30));   //: @(633,160) /sn:0 /w:[ 1 1 0 ] /dr:0
  tran g8(.Z(w9), .I(w4[20:16]));   //: @(296,512) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:0
  MEM g3 (.memWrite(w40), .Address(w23), .write_data(w15), .MemRead(w37), .read_data(w28));   //: @(1165, 137) /sz:(128, 174) /sn:0 /p:[ Ti0>1 Li0>5 Li1>3 Bi0>1 Ro0<0 ]
  //: joint g16 (w25) @(717, 433) /w:[ 1 2 -1 4 ]
  //: joint g17 (w3) @(827, 177) /w:[ 4 6 -1 3 ]
  //: switch g26 (w0) @(-249,690) /sn:0 /w:[ 0 ] /st:0
  EXE g2 (.ALU_operation(w45), .data_read_2(w31), .data_read_1(w16), .PCNext(w3), .INM32(w25), .Zero_signal(w24), .ALU_result(w23), .branch_target(w22));   //: @(867, 86) /sz:(185, 314) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Li2>5 Li3>3 Ro0<0 Ro1<0 Ro2<0 ]
  and g23 (.I0(w36), .I1(w24), .Z(w18));   //: @(1076,59) /sn:0 /w:[ 1 1 0 ]
  READ g1 (.RegWrite(w42), .Read_register_1(w10), .Read_register_2(w9), .Write_register(w8), .mux_RegDst(w11), .Sign_ext_in(w6), .clk(w13), .clr(w0), .Write_data(w32), .Read_data_1(w16), .Read_data_2(w15), .Sign_ext_out(w25));   //: @(404, 335) /sz:(255, 283) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Li2>0 Li3>1 Li4>0 Bi0>0 Bi1>1 Bi2>1 Ro0<0 Ro1<0 Ro2<5 ]
  clock g24 (.Z(w13));   //: @(-253,463) /sn:0 /w:[ 5 ] /omega:100 /phi:0 /duty:50
  mux g18 (.I0(w33), .I1(w30), .S(w14), .Z(w35));   //: @(1210,-62) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:0 /do:0
  tran g10(.Z(w6), .I(w4[15:0]));   //: @(301,571) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  //: joint g25 (w13) @(-146, 463) /w:[ 2 -1 4 1 ]
  tran g6(.Z(w29), .I(w4[25:0]));   //: @(232,429) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:0
  tran g7(.Z(w10), .I(w4[25:21]));   //: @(250,518) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:0
  tran g9(.Z(w8), .I(w4[15:11]));   //: @(344,505) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:0
  tran g22(.Z(w2), .I(w4[31:26]));   //: @(143,482) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:0
  //: joint g12 (w15) @(787, 497) /w:[ 2 4 1 -1 ]
  tran g5(.Z(w19), .I(w3[31:28]));   //: @(546,187) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  mux g11 (.I0(w15), .I1(w25), .S(w41), .Z(w31));   //: @(833,443) /sn:0 /R:1 /w:[ 5 0 1 0 ] /ss:0 /do:0
  //: joint g14 (w23) @(1116, 232) /w:[ 2 4 -1 1 ]
  ctrl g19 (.instruction(w2), .RegWrite(w42), .ALUSrc(w41), .MemWrite(w40), .MemtoReg(w39), .ALUOp(w44), .MemRead(w37), .Branch(w36), .Jump(w14), .RegDst(w11));   //: @(256, -90) /sz:(171, 204) /sn:0 /p:[ Li0>0 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<1 Ro5<0 Ro6<0 Ro7<0 Ro8<0 ]
  tran g21(.Z(w43), .I(w4[5:0]));   //: @(184,427) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:0
  ALUCtrl g20 (.ALUOp(w44), .funct(w43), .ALUCtrl(w45));   //: @(681, -267) /sz:(134, 106) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  mux g15 (.I0(w3), .I1(w22), .S(w18), .Z(w33));   //: @(1122,-42) /sn:0 /R:1 /w:[ 7 1 1 0 ] /ss:0 /do:0
  fetch g0 (.PCNew(w35), .reset(w1), .clk(w13), .Inst(w4), .PCNext(w3));   //: @(-62, 217) /sz:(139, 319) /sn:0 /p:[ Li0>1 Li1>0 Li2>3 Ro0<0 Ro1<0 ]
  mux g13 (.I0(w23), .I1(w28), .S(w39), .Z(w32));   //: @(1378,219) /sn:0 /R:1 /w:[ 3 1 1 0 ] /ss:0 /do:0

endmodule
